module cache_map();



endmodule
